module Sign_Extend
(
	input		[15:0]	Imm,
	
	output	[31:0]	Sign_Ext_Imm
);

	assign Sign_Ext_Imm = {{16{Imm[15]}},Imm};
		
endmodule
