module Decoder
(
	input			[4:0]		Write_Register,
	
	output reg	[31:0]	one_hot
);
	
	always@(*) begin
		case (Write_Register)
			0	:	one_hot = 32'b00000000_00000000_00000000_00000001;
			1	:	one_hot = 32'b00000000_00000000_00000000_00000010;
			2	:	one_hot = 32'b00000000_00000000_00000000_00000100;
			3	:	one_hot = 32'b00000000_00000000_00000000_00001000;
			4	:	one_hot = 32'b00000000_00000000_00000000_00010000;
			5	:	one_hot = 32'b00000000_00000000_00000000_00100000;
			6	:	one_hot = 32'b00000000_00000000_00000000_01000000;
			7	:	one_hot = 32'b00000000_00000000_00000000_10000000;
			8	:	one_hot = 32'b00000000_00000000_00000001_00000000;
			9	:	one_hot = 32'b00000000_00000000_00000010_00000000;
			10	:	one_hot = 32'b00000000_00000000_00000100_00000000;
			11	:	one_hot = 32'b00000000_00000000_00001000_00000000;
			12	:	one_hot = 32'b00000000_00000000_00010000_00000000;
			13	:	one_hot = 32'b00000000_00000000_00100000_00000000;
			14	:	one_hot = 32'b00000000_00000000_01000000_00000000;
			15	:	one_hot = 32'b00000000_00000000_10000000_00000000;
			16	:	one_hot = 32'b00000000_00000001_00000000_00000000;
			17	:	one_hot = 32'b00000000_00000010_00000000_00000000;
			18	:	one_hot = 32'b00000000_00000100_00000000_00000000;
			19	:	one_hot = 32'b00000000_00001000_00000000_00000000;
			20	:	one_hot = 32'b00000000_00010000_00000000_00000000;
			21	:	one_hot = 32'b00000000_00100000_00000000_00000000;
			22	:	one_hot = 32'b00000000_01000000_00000000_00000000;
			23	:	one_hot = 32'b00000000_10000000_00000000_00000000;
			24	:	one_hot = 32'b00000001_00000000_00000000_00000000;
			25	:	one_hot = 32'b00000010_00000000_00000000_00000000;
			26	:	one_hot = 32'b00000100_00000000_00000000_00000000;
			27	:	one_hot = 32'b00001000_00000000_00000000_00000000;
			28	:	one_hot = 32'b00010000_00000000_00000000_00000000;
			29	:	one_hot = 32'b00100000_00000000_00000000_00000000;
			30	:	one_hot = 32'b01000000_00000000_00000000_00000000;
			31	:	one_hot = 32'b10000000_00000000_00000000_00000000;
		endcase
	end	
endmodule
